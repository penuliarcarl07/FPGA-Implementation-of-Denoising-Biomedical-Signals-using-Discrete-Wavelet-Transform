library verilog;
use verilog.vl_types.all;
entity DWT_Algo_tb is
end DWT_Algo_tb;
