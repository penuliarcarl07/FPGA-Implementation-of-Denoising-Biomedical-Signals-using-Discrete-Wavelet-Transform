library verilog;
use verilog.vl_types.all;
entity DWT_db2_3level_tb is
end DWT_db2_3level_tb;
